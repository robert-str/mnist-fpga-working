/*
================================================================================
Isolated Testbench for 2-Hidden-Layer Inference Module
================================================================================

Purpose: Test inference.v in isolation using exact same data preparation as
         Python simulation to eliminate all other error sources.

Model Architecture:
  - Input:  784 pixels (28x28 image, 8-bit signed)
  - Layer 1: 784 → 16 neurons (ReLU activation, right-shift by 7)
  - Layer 2: 16 → 16 neurons (ReLU activation, right-shift by 7)
  - Layer 3: 16 → 10 outputs (no ReLU, no shift)

Strategy:
  1. Load actual weights and biases from .mem files (all 6 BRAMs)
  2. Load preprocessed test vectors generated by Python
  3. Run inference on each test case
  4. Compare results with expected scores from Python simulation
  5. Report any mismatches

Memory Layout:
  - L1 Weights: 12544 bytes (16 neurons × 784 inputs)
  - L1 Biases:  16 × 32-bit
  - L2 Weights: 256 bytes (16 neurons × 16 inputs)
  - L2 Biases:  16 × 32-bit
  - L3 Weights: 160 bytes (10 classes × 16 inputs)
  - L3 Biases:  10 × 32-bit

================================================================================
*/

`timescale 1ns / 1ps

module tb_inference();

    // Parameters
    parameter NUM_PIXELS = 784;
    parameter L1_NEURONS = 16;
    parameter L2_NEURONS = 16;
    parameter NUM_CLASSES = 10;
    parameter NUM_TEST_CASES = 100;
    
    // Clock and Reset
    reg clk;
    reg rst;
    
    // Layer 1 Memory Interfaces
    wire [13:0] L1_weight_addr;
    reg  [7:0]  L1_weight_data;
    wire [3:0]  L1_bias_addr;
    reg  [31:0] L1_bias_data;
    
    // Layer 2 Memory Interfaces
    wire [7:0]  L2_weight_addr;
    reg  [7:0]  L2_weight_data;
    wire [3:0]  L2_bias_addr;
    reg  [31:0] L2_bias_data;
    
    // Layer 3 Memory Interfaces
    wire [7:0]  L3_weight_addr;
    reg  [7:0]  L3_weight_data;
    wire [3:0]  L3_bias_addr;
    reg  [31:0] L3_bias_data;
    
    // Input Image Interface
    wire [9:0]  input_addr;
    reg  [7:0]  input_pixel;
    
    // Control
    reg weights_ready;
    reg start_inference;
    
    // Outputs
    wire [3:0] predicted_digit;
    wire inference_done;
    wire busy;
    
    // Class scores
    wire signed [31:0] class_score_0;
    wire signed [31:0] class_score_1;
    wire signed [31:0] class_score_2;
    wire signed [31:0] class_score_3;
    wire signed [31:0] class_score_4;
    wire signed [31:0] class_score_5;
    wire signed [31:0] class_score_6;
    wire signed [31:0] class_score_7;
    wire signed [31:0] class_score_8;
    wire signed [31:0] class_score_9;
    
    // ========================================================================
    // Memory Storage
    // ========================================================================
    
    // Weight and Bias memories
    reg [7:0]  L1_weights_mem [0:12543];   // 16 × 784 = 12544
    reg [31:0] L1_biases_mem  [0:15];      // 16 biases
    reg [7:0]  L2_weights_mem [0:255];     // 16 × 16 = 256
    reg [31:0] L2_biases_mem  [0:15];      // 16 biases
    reg [7:0]  L3_weights_mem [0:159];     // 10 × 16 = 160
    reg [31:0] L3_biases_mem  [0:9];       // 10 biases
    
    // Test vector storage (flattened for $readmemh)
    reg [7:0] test_pixels_flat [0:78399];           // 100 tests × 784 pixels
    reg signed [31:0] expected_scores_flat [0:999]; // 100 tests × 10 scores
    reg [3:0] expected_predictions [0:99];
    reg [3:0] true_labels [0:99];
    
    // Test control
    integer test_idx;
    integer pass_count;
    integer fail_count;
    integer pred_match_count;
    integer j;
    integer file_check;
    reg signed [31:0] max_error;
    reg scores_match;
    reg signed [31:0] fpga_scores [0:9];
    reg signed [31:0] diff;
    
    // ========================================================================
    // Instantiate the Unit Under Test (UUT)
    // ========================================================================
    inference uut (
        .clk(clk),
        .rst(rst),
        
        // Layer 1 interface
        .L1_weight_addr(L1_weight_addr),
        .L1_weight_data(L1_weight_data),
        .L1_bias_addr(L1_bias_addr),
        .L1_bias_data(L1_bias_data),
        
        // Layer 2 interface
        .L2_weight_addr(L2_weight_addr),
        .L2_weight_data(L2_weight_data),
        .L2_bias_addr(L2_bias_addr),
        .L2_bias_data(L2_bias_data),
        
        // Layer 3 interface
        .L3_weight_addr(L3_weight_addr),
        .L3_weight_data(L3_weight_data),
        .L3_bias_addr(L3_bias_addr),
        .L3_bias_data(L3_bias_data),
        
        // Control
        .weights_ready(weights_ready),
        .start_inference(start_inference),
        .input_pixel(input_pixel),
        .input_addr(input_addr),
        
        // Outputs
        .predicted_digit(predicted_digit),
        .inference_done(inference_done),
        .busy(busy),
        
        // Class scores
        .class_score_0(class_score_0),
        .class_score_1(class_score_1),
        .class_score_2(class_score_2),
        .class_score_3(class_score_3),
        .class_score_4(class_score_4),
        .class_score_5(class_score_5),
        .class_score_6(class_score_6),
        .class_score_7(class_score_7),
        .class_score_8(class_score_8),
        .class_score_9(class_score_9)
    );
    
    // Clock Generation: 100MHz (10ns period)
    always #5 clk = ~clk;
    
    // ========================================================================
    // Memory Interface Logic - Simulates BRAM behavior with 1-cycle latency
    // ========================================================================
    
    // Layer 1 Weight Memory
    always @(posedge clk) begin
        if (L1_weight_addr < 12544)
            L1_weight_data <= L1_weights_mem[L1_weight_addr];
        else
            L1_weight_data <= 8'd0;
    end
    
    // Layer 1 Bias Memory
    always @(posedge clk) begin
        if (L1_bias_addr < 16)
            L1_bias_data <= L1_biases_mem[L1_bias_addr];
        else
            L1_bias_data <= 32'd0;
    end
    
    // Layer 2 Weight Memory
    always @(posedge clk) begin
        if (L2_weight_addr < 256)
            L2_weight_data <= L2_weights_mem[L2_weight_addr];
        else
            L2_weight_data <= 8'd0;
    end
    
    // Layer 2 Bias Memory
    always @(posedge clk) begin
        if (L2_bias_addr < 16)
            L2_bias_data <= L2_biases_mem[L2_bias_addr];
        else
            L2_bias_data <= 32'd0;
    end
    
    // Layer 3 Weight Memory
    always @(posedge clk) begin
        if (L3_weight_addr < 160)
            L3_weight_data <= L3_weights_mem[L3_weight_addr];
        else
            L3_weight_data <= 8'd0;
    end
    
    // Layer 3 Bias Memory
    always @(posedge clk) begin
        if (L3_bias_addr < 10)
            L3_bias_data <= L3_biases_mem[L3_bias_addr];
        else
            L3_bias_data <= 32'd0;
    end
    
    // Input Pixel Memory (access flattened array based on current test)
    always @(posedge clk) begin
        if (input_addr < 784)
            input_pixel <= test_pixels_flat[test_idx * 784 + input_addr];
        else
            input_pixel <= 8'd0;
    end
    
    // ========================================================================
    // Load Memory Files
    // ========================================================================
    initial begin
        $display("================================================================================");
        $display("Loading Memory Files...");
        $display("================================================================================");
        $display("Current working directory for file loading:");
        $display("  (Vivado runs from simulation directory)");
        $display("");
        
        // Load L1 weights with error checking
        file_check = $fopen("L1_weights.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open L1_weights.mem");
            $display("  Make sure L1_weights.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("L1_weights.mem", L1_weights_mem);
        $display("  [OK] Loaded L1 weights: 12544 entries");
        
        // Load L1 biases with error checking
        file_check = $fopen("L1_biases.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open L1_biases.mem");
            $display("  Make sure L1_biases.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("L1_biases.mem", L1_biases_mem);
        $display("  [OK] Loaded L1 biases: 16 entries");
        
        // Load L2 weights with error checking
        file_check = $fopen("L2_weights.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open L2_weights.mem");
            $display("  Make sure L2_weights.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("L2_weights.mem", L2_weights_mem);
        $display("  [OK] Loaded L2 weights: 256 entries");
        
        // Load L2 biases with error checking
        file_check = $fopen("L2_biases.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open L2_biases.mem");
            $display("  Make sure L2_biases.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("L2_biases.mem", L2_biases_mem);
        $display("  [OK] Loaded L2 biases: 16 entries");
        
        // Load L3 weights with error checking
        file_check = $fopen("L3_weights.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open L3_weights.mem");
            $display("  Make sure L3_weights.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("L3_weights.mem", L3_weights_mem);
        $display("  [OK] Loaded L3 weights: 160 entries");
        
        // Load L3 biases with error checking
        file_check = $fopen("L3_biases.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open L3_biases.mem");
            $display("  Make sure L3_biases.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("L3_biases.mem", L3_biases_mem);
        $display("  [OK] Loaded L3 biases: 10 entries");
        
        // Load test vectors (flattened format) with error checking
        file_check = $fopen("test_vectors_pixels.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_pixels.mem");
            $display("  Make sure test_vectors_pixels.mem is added as simulation source");
            $display("  Run generate_test_vectors.py first!");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_pixels.mem", test_pixels_flat);
        $display("  [OK] Loaded pixel vectors: 78400 values");
        
        file_check = $fopen("test_vectors_scores.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_scores.mem");
            $display("  Make sure test_vectors_scores.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_scores.mem", expected_scores_flat);
        $display("  [OK] Loaded score vectors: 1000 values");
        
        file_check = $fopen("test_vectors_meta.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_meta.mem");
            $display("  Make sure test_vectors_meta.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_meta.mem", expected_predictions);
        $display("  [OK] Loaded predictions: 100 values");
        
        file_check = $fopen("test_vectors_labels.mem", "r");
        if (file_check == 0) begin
            $display("ERROR: Cannot open test_vectors_labels.mem");
            $display("  Make sure test_vectors_labels.mem is added as simulation source");
            $finish;
        end
        $fclose(file_check);
        $readmemh("test_vectors_labels.mem", true_labels);
        $display("  [OK] Loaded labels: 100 values");
        
        $display("  [OK] Loaded test vectors: %0d test cases", NUM_TEST_CASES);
        
        $display("================================================================================\n");
    end
    
    // ========================================================================
    // Test Sequence
    // ========================================================================
    initial begin
        $display("================================================================================");
        $display("Isolated Testbench for 2-Hidden-Layer inference.v");
        $display("================================================================================");
        $display("Testing inference.v in complete isolation using:");
        $display("  - Real weight and bias files from training (L1, L2, L3)");
        $display("  - Preprocessed test vectors from Python (same as UART sends)");
        $display("  - Expected scores from Python simulation");
        $display("================================================================================\n");
        
        // Initialize
        clk = 0;
        rst = 1;
        weights_ready = 0;
        start_inference = 0;
        test_idx = 0;
        pass_count = 0;
        fail_count = 0;
        pred_match_count = 0;
        
        // Reset
        #100;
        rst = 0;
        #20;
        
        $display("[%0t] Starting Isolated Inference Tests\n", $time);
        weights_ready = 1;
        
        // Run tests on all test cases
        for (test_idx = 0; test_idx < NUM_TEST_CASES; test_idx = test_idx + 1) begin
            $display("================================================================================");
            $display("Test Case %0d / %0d", test_idx + 1, NUM_TEST_CASES);
            $display("================================================================================");
            $display("  True Label:         %0d", true_labels[test_idx]);
            $display("  Expected Pred:      %0d (from Python sim)", expected_predictions[test_idx]);
            
            // Start inference
            #10 start_inference = 1;
            #10 start_inference = 0;
            
            // Wait for completion
            wait(inference_done);
            #20;
            
            // Collect FPGA scores
            fpga_scores[0] = class_score_0;
            fpga_scores[1] = class_score_1;
            fpga_scores[2] = class_score_2;
            fpga_scores[3] = class_score_3;
            fpga_scores[4] = class_score_4;
            fpga_scores[5] = class_score_5;
            fpga_scores[6] = class_score_6;
            fpga_scores[7] = class_score_7;
            fpga_scores[8] = class_score_8;
            fpga_scores[9] = class_score_9;
            
            // Verify results
            $display("  FPGA Pred:          %0d", predicted_digit);
            $display("\n  Score Comparison:");
            $display("  Class | Expected      | FPGA          | Difference");
            $display("  ------|---------------|---------------|---------------");
            
            scores_match = 1;
            max_error = 0;
            
            // Compare all class scores
            for (j = 0; j < 10; j = j + 1) begin
                diff = fpga_scores[j] - expected_scores_flat[test_idx * 10 + j];
                
                if (fpga_scores[j] !== expected_scores_flat[test_idx * 10 + j]) begin
                    scores_match = 0;
                    if ($signed(diff) < 0) begin
                        if (-diff > max_error) max_error = -diff;
                    end else begin
                        if (diff > max_error) max_error = diff;
                    end
                end
                
                $display("    %0d   | %13d | %13d | %13d %s",
                        j, expected_scores_flat[test_idx * 10 + j], fpga_scores[j], diff,
                        (fpga_scores[j] !== expected_scores_flat[test_idx * 10 + j]) ? "<-- MISMATCH" : "");
            end
            
            // Track prediction match separately
            if (predicted_digit == expected_predictions[test_idx]) begin
                pred_match_count = pred_match_count + 1;
            end
            
            // Check overall result
            $display("\n  Max Score Error:    %0d", max_error);
            $display("  Scores Match:       %s", scores_match ? "YES" : "NO");
            $display("  Pred Match:         %s", (predicted_digit == expected_predictions[test_idx]) ? "YES" : "NO");
            
            if (scores_match && (predicted_digit == expected_predictions[test_idx])) begin
                $display("  Result:             PASS");
                pass_count = pass_count + 1;
            end else begin
                $display("  Result:             FAIL");
                fail_count = fail_count + 1;
            end
            
            $display("");
            
            // Small delay between tests
            #50;
        end
        
        // Final Summary
        $display("\n================================================================================");
        $display("FINAL RESULTS");
        $display("================================================================================");
        $display("Total Tests:             %0d", NUM_TEST_CASES);
        $display("Exact Score Matches:     %0d", pass_count);
        $display("Score Mismatches:        %0d", fail_count);
        $display("Prediction Matches:      %0d (%.1f%%)", pred_match_count, (pred_match_count * 100.0) / NUM_TEST_CASES);
        $display("================================================================================");
        
        if (fail_count == 0) begin
            $display("\nALL TESTS PASSED - EXACT SCORE MATCH");
            $display("inference.v is computing correctly!");
            $display("The mismatch problem is NOT in inference.v");
            $display("Check other modules: UART, image_loader, weight_loader, etc.");
        end else if (pred_match_count == NUM_TEST_CASES) begin
            $display("\nPREDICTION MATCH BUT SCORE DIFFERENCES");
            $display("The predictions are correct but scores differ slightly.");
            $display("This may be due to minor numerical differences that don't affect the result.");
        end else begin
            $display("\nTESTS FAILED");
            $display("inference.v has computation errors!");
            $display("Review the detailed comparisons above.");
            $display("Possible issues:");
            $display("  - Pipeline timing bug");
            $display("  - Sign extension error");
            $display("  - Accumulator overflow handling");
            $display("  - Weight/bias memory addressing");
            $display("  - Right-shift implementation");
        end
        $display("================================================================================\n");
        
        #100;
        $finish;
    end
    
    // Timeout watchdog
    initial begin
        #500000000;  // 500ms timeout (3-layer network takes longer)
        $display("\nERROR: Simulation timeout!");
        $finish;
    end

endmodule


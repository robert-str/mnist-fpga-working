module image_loader (
    input wire clk,
    input wire rst,
    input wire weights_loaded,
    input wire [7:0] rx_data,
    input wire rx_ready,
    output reg [9:0] wr_addr,
    output reg [7:0] wr_data,
    output reg wr_en,
    output reg image_loaded
);
    localparam IMG_END1 = 8'h66;
    localparam IMG_END2 = 8'hBB;
    localparam IMG_SIZE = 784;

    localparam STATE_RECEIVING = 2'd0;
    localparam STATE_DONE      = 2'd1;

    reg [1:0] state;
    reg [9:0] byte_count;
    reg [7:0] prev_byte;

    // === NEW: Input Registration Logic ===
    // This captures the wire inputs into registers to fix timing/glitches
    reg [7:0] rx_data_reg;
    reg rx_ready_reg;

    always @(posedge clk) begin
        rx_data_reg <= rx_data;
        rx_ready_reg <= rx_ready;
    end
    // ======================================

    always @(posedge clk) begin
        if (rst) begin
            state <= STATE_RECEIVING;
            wr_addr <= 0;
            wr_data <= 0;
            wr_en <= 0;
            byte_count <= 0;
            prev_byte <= 0;
            image_loaded <= 0;
        end else begin
            wr_en <= 0;
            image_loaded <= 0;
            
            if (weights_loaded) begin
                case (state)
                    STATE_RECEIVING: begin
                        // CHANGE: Use the REGISTERED signal (rx_ready_reg)
                        if (rx_ready_reg) begin
                            // 1. Write previous byte (if exists)
                            if (byte_count > 0 && byte_count <= IMG_SIZE) begin
                                wr_addr <= byte_count - 1;
                                wr_data <= prev_byte;
                                wr_en <= 1;
                            end
                            
                            // 2. Check End Condition (Use registered data)
                            // Note: We check rx_data_reg here!
                            if (byte_count >= IMG_SIZE && prev_byte == IMG_END1 && rx_data_reg == IMG_END2) begin
                                state <= STATE_DONE;
                                image_loaded <= 1;
                                // DEBUG PRINT
                                $display("[%t] IMAGE LOADED SUCCESS! Count: %d", $time, byte_count);
                            end else begin
                                // 3. Pipeline current byte
                                byte_count <= byte_count + 1;
                                prev_byte <= rx_data_reg;
                            end
                        end
                    end
                    
                    STATE_DONE: begin
                        state <= STATE_RECEIVING;
                        byte_count <= 0;
                        prev_byte <= 0;
                    end
                endcase
            end
        end
    end
endmodule
